`include "rom32x4.v"

`default_nettype none

module romhw (
  input wire clk,
  output wire [7:0] leds
);

localparam ADDR = 5'h5;

rom32x4
  ROM (.clk(clk), .addr(ADDR), .data(leds[3:0]));

assign leds[7:4] = 0;

endmodule
